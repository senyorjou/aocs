module main

fn main() {
	println('Advent of Code 2025 - VLang Project')
	println('Run specific day solutions using `v run src/dayXX.v`')
}

